class







endclass
