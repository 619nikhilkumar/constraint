class



function
  endfunction



endclass
